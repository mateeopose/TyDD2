library verilog;
use verilog.vl_types.all;
entity multi2consigno_vlg_vec_tst is
end multi2consigno_vlg_vec_tst;
