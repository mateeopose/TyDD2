library verilog;
use verilog.vl_types.all;
entity circuitoi2c_vlg_vec_tst is
end circuitoi2c_vlg_vec_tst;
