library verilog;
use verilog.vl_types.all;
entity Sumador_Completo_vlg_vec_tst is
end Sumador_Completo_vlg_vec_tst;
