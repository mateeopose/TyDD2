library verilog;
use verilog.vl_types.all;
entity comparador_vlg_check_tst is
    port(
        soy             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end comparador_vlg_check_tst;
