-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Oct 26 18:33:55 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY i2c IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        sda : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        hab_dir : OUT STD_LOGIC;
        hab_dat : OUT STD_LOGIC;
        ackout : OUT STD_LOGIC
    );
END i2c;

ARCHITECTURE BEHAVIOR OF i2c IS
    TYPE type_fstate IS (Idle,guarda_direc,RW,ACK,guarda_dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= Idle;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,sda,fin_dir,soy,fin_dato)
    BEGIN
        hab_dir <= '0';
        hab_dat <= '0';
        ackout <= '0';
        CASE fstate IS
            WHEN Idle =>
                IF ((sda = '0')) THEN
                    reg_fstate <= guarda_direc;
                ELSIF ((sda = '1')) THEN
                    reg_fstate <= Idle;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Idle;
                END IF;
            WHEN guarda_direc =>
                IF ((fin_dir = '0')) THEN
                    reg_fstate <= guarda_direc;
                ELSIF (((fin_dir = '1') AND (soy = '0'))) THEN
                    reg_fstate <= Idle;
                ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                    reg_fstate <= RW;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= guarda_direc;
                END IF;

                hab_dir <= '1';
            WHEN RW =>
                reg_fstate <= ACK;
            WHEN ACK =>
                reg_fstate <= guarda_dato;

                ackout <= '1';
            WHEN guarda_dato =>
                IF ((fin_dato = '0')) THEN
                    reg_fstate <= guarda_dato;
                ELSIF ((fin_dato = '1')) THEN
                    reg_fstate <= Idle;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= guarda_dato;
                END IF;

                hab_dat <= '1';
            WHEN OTHERS => 
                hab_dir <= 'X';
                hab_dat <= 'X';
                ackout <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
