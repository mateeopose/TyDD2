library verilog;
use verilog.vl_types.all;
entity multi2sinsigno_vlg_vec_tst is
end multi2sinsigno_vlg_vec_tst;
