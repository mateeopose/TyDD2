library verilog;
use verilog.vl_types.all;
entity multi2sinsigno_vlg_check_tst is
    port(
        Out0            : in     vl_logic;
        Out1            : in     vl_logic;
        Out2            : in     vl_logic;
        Out3            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end multi2sinsigno_vlg_check_tst;
