-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Thu Oct 30 14:58:20 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY multi2consigno IS 
	PORT
	(
		b0 :  IN  STD_LOGIC;
		a0 :  IN  STD_LOGIC;
		Cin :  IN  STD_LOGIC;
		b1 :  IN  STD_LOGIC;
		a1 :  IN  STD_LOGIC;
		PRN :  IN  STD_LOGIC;
		CLRN :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		Out0 :  OUT  STD_LOGIC;
		Out1 :  OUT  STD_LOGIC;
		Out3 :  OUT  STD_LOGIC;
		Out2 :  OUT  STD_LOGIC;
		prueba :  OUT  STD_LOGIC
	);
END multi2consigno;

ARCHITECTURE bdf_type OF multi2consigno IS 

COMPONENT sumador_completo
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 Cout : OUT STD_LOGIC;
		 Sum : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;


BEGIN 
prueba <= SYNTHESIZED_WIRE_18;
SYNTHESIZED_WIRE_20 <= '1';



PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	SYNTHESIZED_WIRE_21 <= '0';
ELSIF (PRN = '0') THEN
	SYNTHESIZED_WIRE_21 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_21 <= a0;
END IF;
END PROCESS;



PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	SYNTHESIZED_WIRE_24 <= '0';
ELSIF (PRN = '0') THEN
	SYNTHESIZED_WIRE_24 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_24 <= b1;
END IF;
END PROCESS;


PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	SYNTHESIZED_WIRE_22 <= '0';
ELSIF (PRN = '0') THEN
	SYNTHESIZED_WIRE_22 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_22 <= a1;
END IF;
END PROCESS;


PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	Out0 <= '0';
ELSIF (PRN = '0') THEN
	Out0 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	Out0 <= SYNTHESIZED_WIRE_0;
END IF;
END PROCESS;


PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	Out1 <= '0';
ELSIF (PRN = '0') THEN
	Out1 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	Out1 <= SYNTHESIZED_WIRE_1;
END IF;
END PROCESS;


PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	Out2 <= '0';
ELSIF (PRN = '0') THEN
	Out2 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	Out2 <= SYNTHESIZED_WIRE_2;
END IF;
END PROCESS;


PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	Out3 <= '0';
ELSIF (PRN = '0') THEN
	Out3 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	Out3 <= SYNTHESIZED_WIRE_3;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_19 <= NOT(SYNTHESIZED_WIRE_21);



SYNTHESIZED_WIRE_23 <= NOT(SYNTHESIZED_WIRE_22);



b2v_inst18 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_4,
		 B => SYNTHESIZED_WIRE_23,
		 Sum => SYNTHESIZED_WIRE_9,
		 Cin => '0',
		 cout => open );


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_24;


b2v_inst2 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_25,
		 B => SYNTHESIZED_WIRE_8,
		 Cin => Cin,
		 Cout => SYNTHESIZED_WIRE_16,
		 Sum => SYNTHESIZED_WIRE_1);


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_9 AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_24 AND SYNTHESIZED_WIRE_23;


b2v_inst22 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_25,
		 B => SYNTHESIZED_WIRE_12,
		 Cin => SYNTHESIZED_WIRE_13,
		 Sum => SYNTHESIZED_WIRE_17);


b2v_inst3 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_25,
		 B => SYNTHESIZED_WIRE_15,
		 Cin => SYNTHESIZED_WIRE_16,
		 Cout => SYNTHESIZED_WIRE_13,
		 Sum => SYNTHESIZED_WIRE_2);


SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_17 AND SYNTHESIZED_WIRE_18;


b2v_inst8 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_19,
		 B => SYNTHESIZED_WIRE_20,
		 Cin => Cin,
		 Cout => SYNTHESIZED_WIRE_4,
		 Sum => SYNTHESIZED_WIRE_6);


PROCESS(CLK,CLRN,PRN)
BEGIN
IF (CLRN = '0') THEN
	SYNTHESIZED_WIRE_26 <= '0';
ELSIF (PRN = '0') THEN
	SYNTHESIZED_WIRE_26 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_26 <= b0;
END IF;
END PROCESS;


END bdf_type;