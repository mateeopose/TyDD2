library verilog;
use verilog.vl_types.all;
entity Multimodca2_vlg_vec_tst is
end Multimodca2_vlg_vec_tst;
