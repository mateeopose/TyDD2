library verilog;
use verilog.vl_types.all;
entity i2c_vlg_vec_tst is
end i2c_vlg_vec_tst;
