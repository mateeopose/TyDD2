library ieee;
use ieee.std_logic_1164.all;

entity Sumador_Completo is
	port( A: in std_logic;
			B: in std_logic;
			Cin: in std_logic;
			Cout: out std_logic;
			
	