library verilog;
use verilog.vl_types.all;
entity Multimodca2_vlg_sample_tst is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        b0              : in     vl_logic;
        b1              : in     vl_logic;
        Cin             : in     vl_logic;
        CLK             : in     vl_logic;
        CLRN            : in     vl_logic;
        PRN             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Multimodca2_vlg_sample_tst;
