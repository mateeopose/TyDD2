library verilog;
use verilog.vl_types.all;
entity maqestados_vlg_vec_tst is
end maqestados_vlg_vec_tst;
